package counter_pkg;
   `include "tester.svh"
   `include "ctr_checker.svh"
   `include "monitor.svh"
  
endpackage // counter_pkg

